library ieee;

use ieee.std_logic_1164.all;

package xbar_package is
	
end xbar_package;